`timescale 1ns/1ns

module testbench_top;
   reg clk, rst, start;
   reg [9:0] A, B;
   wire ov;
   wire [9:0] Q;
   wire busy , valid,dvz;
   div_top uut (clk,start,A, B, Q, busy, valid,ov,dvz);

   assign clk = 0;
   initial begin forever #5 clk = ~clk; end

   initial
   begin
      // Devide by zero :
      A = 10'b1101010000;
      B = 10'b0;
      rst = 1; start = 0; 
     #10 rst = 0; start = 1;#10 start=0; #380;
      // Main Tests: 
      A = 10'b0000101010;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0110101111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1100000100;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0101110010;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0001000100;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1001110111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0001100011;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0101001111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1011110100;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1001010001;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0000101000;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0110000001;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1010000111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1000011110;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1000101110;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0110111111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1111110011;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0101010111;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0110000111;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0010011100;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0010010100;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111001110;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1011001001;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111000110;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111000110;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1001100111;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1000001011;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1000101101;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0000010110;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1111010010;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1111000010;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1111010111;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111111111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111010101;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1110010001;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1010000001;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1011111110;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1101100101;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1010010101;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0110011000;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0000111101;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0010011011;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1000011000;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0100111011;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1101010110;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0100100001;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0100101111;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0100100110;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1111010001;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1101111110;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0100100111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0000111111;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0000010011;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1000010000;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0000100110;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0110000000;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1111110011;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0000010101;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0000110000;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1000100101;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111100101;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111100101;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1101001000;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1101001110;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111111111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1101110101;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0001100111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0010101101;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1001010011;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0100110000;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1011100000;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1110010101;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0001001010;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1110000000;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1000101111;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0110000100;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1010000100;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1001001000;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1101001010;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0110101100;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111100110;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1101010000;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111011111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111111100;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1111111111;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111010000;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0100001000;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111010110;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1010000110;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1111111110;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1000110100;
      B = 10'b0000010000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0101010010;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1111000000;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0111110101;
      B = 10'b0000011000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0110111111;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b1011110001;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0101111010;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0100010110;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0000111100;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;

      A = 10'b0000010011;
      B = 10'b0000001000;
      rst = 1; start = 0;
      #10 rst = 0; start = 1;#10 start=0; #380;


      $stop;
   end

endmodule
